library ieee;

package instructions_types is

	type instruction_type is (INVALID, DP_R, DP_I, LS, BBL, STP);

end package;